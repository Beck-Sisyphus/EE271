library verilog;
use verilog.vl_types.all;
entity seg7_testbench is
end seg7_testbench;
