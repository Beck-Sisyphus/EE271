library verilog;
use verilog.vl_types.all;
entity adder_testbench is
end adder_testbench;
