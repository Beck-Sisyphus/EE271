// Beck Pang, EE 271 Lab 4
module highLevelDesign (HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, U, P, C);